parameter X = 2;

module top(b);
input b;
parameter Y = 3;
endmodule

