module top(output [17:0] b);
wire a = 100_000.0;
assign b = 123_456.0;
endmodule

