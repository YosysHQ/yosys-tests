module testbench;
    reg clk;

    initial begin
       //  $dumpfile("testbench.vcd");
       //  $dumpvars(0, testbench);

        #5 clk = 0;
        repeat (10000) begin
            #5 clk = 1;
            #5 clk = 0;
        end

        $display("OKAY");
    end


    reg [7:0] data_a = 0;
	reg [7:0] data_b = 0;
	reg [5:0] addr_a = 0;
	reg [5:0] addr_b = 0;
    reg we_a = 0;
	reg we_b = 1;
    reg re_a = 1;
	reg re_b = 1;
	wire [7:0] q_a,q_b;
	reg mem_init = 0;

	reg [7:0] pq_a,pq_b;

    top uut (
    .data_a(data_a),
	.data_b(data_b),
	.addr_a(addr_a),
	.addr_b(addr_b),
	.we_a(we_a),
	.we_b(we_b),
	.re_a(re_a),
	.re_b(re_b),
	.clk(clk),
	.q_a(q_a),
	.q_b(q_b)
    );

    always @(posedge clk) begin
    #3;
    data_a <= data_a + 17;
    data_b <= data_b + 5;

    addr_a <= addr_a + 1;
    addr_b <= addr_b + 1;
    end

    always @(posedge addr_a) begin
    #10;
        if(addr_a > 6'h3E)
            mem_init <= 1;
    end

	always @(posedge clk) begin
    //#3;
    we_a <= !we_a;
    we_b <= !we_b;
    end

    // Declare the RAM variable for check
	reg [7:0] ram[63:0];

	// Port A for check
	always @ (posedge clk)
	begin
		if (we_a)
		begin
			ram[addr_a] <= data_a;
			pq_a <= data_a;
		end
		if (re_b)
		begin
			pq_a <= ram[addr_a];
		end
	end

	// Port B for check
	always @ (posedge clk)
	begin
		if (we_b)
		begin
			ram[addr_b] <= data_b;
			pq_b <= data_b;
		end
		if (re_b)
		begin
			pq_b <= ram[addr_b];
		end
	end

	uut_mem_checker port_a_test(.clk(clk), .init(mem_init), .en(!we_a), .A(q_a), .B(pq_a));
    uut_mem_checker port_b_test(.clk(clk), .init(mem_init), .en(!we_b), .A(q_b), .B(pq_b));

endmodule

module uut_mem_checker(input clk, input init, input en, input [7:0] A, input [7:0] B);
    always @(posedge clk)
    begin
        #1;
        if (en == 1 & init == 1 & A !== B)
        begin
            $display("ERROR: ASSERTION FAILED in %m:",$time," ",A," ",B);
            $stop;
        end
    end
endmodule
