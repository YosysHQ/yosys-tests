`define N 131
