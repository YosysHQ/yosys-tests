module top ;
enum {A, B} x;
endmodule
