module top
(
 input x
 );

endmodule

module top1
(
 input x
 );

endmodule
